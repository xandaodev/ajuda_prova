aqui vai ser o process
